module Pc_a( IM , clk , Reset , )
